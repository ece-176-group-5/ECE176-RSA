library verilog;
use verilog.vl_types.all;
entity RSA_TB is
end RSA_TB;
