library verilog;
use verilog.vl_types.all;
entity RSA_2_tb is
end RSA_2_tb;
