// Subtracts 1 from 2 inputted prime numbers
module Subtractor_2_input(
  output p_sub,
  output q_sub,
  input p,
  input q);
  
  assign p_sub=p-1;
  assign q_sub=q-1;
endmodule
