module Prime_Number_Generator(
  output p,
  output q,
  output e
  );

parameter n;  // Limit for a prime number



endmodule